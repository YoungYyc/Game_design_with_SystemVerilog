///test///

module top_ver (
input    q, p,
output   out, );
bottom_vhdl u1 (.a(q), .b(p), .c(out));

endmodule


